LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY decoder IS
	PORT (
		-- Input ports
		input : IN STD_LOGIC_VECTOR(7 DOWNTO 0);

		-- Output ports
		habilitaDisplay : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		habilitaRam : OUT STD_LOGIC;
		habilitaBaseDeTempo : OUT STD_LOGIC;
		clearBaseDeTempo : OUT STD_LOGIC;
		habilitaButton : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		habilitaSwitches : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE behavior OF decoder IS

BEGIN

	-- Habilita da RAM atrelado ao bit mais significativo do endereço
	habilitaRam <= '1' WHEN input(7) = '1' ELSE
		'0';

	habilitaDisplay <= "000001" WHEN input = "00000000" ELSE --Display 0
		"000010" WHEN input = "00000001" ELSE --Display 1
		"000100" WHEN input = "00000010" ELSE --Display 2
		"001000" WHEN input = "00000011" ELSE --Display 3
		"010000" WHEN input = "00000100" ELSE --Display 4
		"100000" WHEN input = "00000101" ELSE --Display 5
		"000000";

	habilitaBaseDeTempo <= '1' WHEN input = "00000110" ELSE
		'0'; -- habilita base de tempo

	clearBaseDeTempo <= '1' WHEN input = "00000111" ELSE
		'0'; -- clear base de tempo

	habilitaButton <= "0001" WHEN input = "00001000" ELSE -- Button 3 
		"0010" WHEN input = "00001001" ELSE -- Button 2
		"0100" WHEN input = "00001010" ELSE -- Button 1
		"1000" WHEN input = "00001011" ELSE -- Button 0
		"0000";
		
	habilitaSwitches <= "000000001" WHEN input = "00001100" ELSE -- Switch 0
		"000000010" WHEN input = "00001101" ELSE -- Switch 1
		"000000100" WHEN input = "00001110" ELSE -- Switch 2
		"000001000" WHEN input = "00001111" ELSE -- Switch 3
		"000010000" WHEN input = "00010000" ELSE -- Switch 4
		"000100000" WHEN input = "00010001" ELSE -- Switch 5
		"001000000" WHEN input = "00010010" ELSE -- Switch 6
		"010000000" WHEN input = "00010011" ELSE -- Switch 7
		"100000000" WHEN input = "00010100" ELSE -- Switch 8
		"000000000";

END ARCHITECTURE;